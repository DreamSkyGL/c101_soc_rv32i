//-----------------------------------------------------------------------------
//   Copyright 2022 GanLing, 1577959692@qq.com
//
//   Licensed under the Apache License, Version 2.0 (the "License");
//   you may not use this file except in compliance with the License.
//   You may obtain a copy of the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in writing, software
//   distributed under the License is distributed on an "AS IS" BASIS,
//   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
//   See the License for the specific language governing permissions and
//   limitations under the License.
//-----------------------------------------------------------------------------

module rst_n_sync(
  input   clk,
  input   rst_n_async,
  output  rst_n_sync
);

reg   r1;
reg   r2;

always @ (posedge clk or negedge rst_n_async) begin
  if(!rst_n_async) begin
    r1  <=  1'b0;
    r2  <=  1'b0;
  end
  else begin
    r1  <=  1'b1;
    r2  <=  r1;
  end
end

assign  rst_n_sync  = r2;

endmodule

